A|B|C|D|E|F
1|2||-10|5|6
|8|9|10||12
13|14||16|17|18
-5||15|55|120|
20|39||41|101|90
25||100||22|77
